<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,0,122.4,-60.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>28.5,-3.5</position>
<gparam>LABEL_TEXT Full Adder Using Nand Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>BA_NAND2</type>
<position>17,-23</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>31.5,-13</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>30,-31.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND2</type>
<position>41.5,-22.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>60.5,-12.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND2</type>
<position>61,-32</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND2</type>
<position>50.5,-22.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>BA_NAND2</type>
<position>70.5,-22.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>8,-18.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>8,-27.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>16.5,-40.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_NAND2</type>
<position>65,-41.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>69,-41.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>74.5,-22.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_LABEL</type>
<position>5.5,-18</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_LABEL</type>
<position>5.5,-27</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>11,-40</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>80,-22</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>74.5,-41</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-32.5,14,-24</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-32.5 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-27.5,14,-27.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-32.5,27,-32.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-22,14,-12</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-18.5,14,-18.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-12,28.5,-12</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-21.5,36.5,-13</points>
<intersection>-21.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-21.5,38.5,-21.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-13,36.5,-13</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-31.5,35.5,-23.5</points>
<intersection>-31.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-31.5,35.5,-31.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-23.5,38.5,-23.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-22.5,46,-21.5</points>
<intersection>-22.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-22.5,46,-22.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-21.5,47.5,-21.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,-21.5,47.5,-11.5</points>
<intersection>-21.5 2</intersection>
<intersection>-11.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-11.5,57.5,-11.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>47.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-40.5,46,-23.5</points>
<intersection>-40.5 1</intersection>
<intersection>-33 3</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-40.5,46,-40.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-23.5,47.5,-23.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>46,-33,58,-33</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-42.5,24.5,-14</points>
<intersection>-42.5 5</intersection>
<intersection>-30.5 1</intersection>
<intersection>-23 2</intersection>
<intersection>-14 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-30.5,27,-30.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-23,24.5,-23</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>24.5,-42.5,62,-42.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>24.5,-14,28.5,-14</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-40.5,56,-13.5</points>
<intersection>-40.5 1</intersection>
<intersection>-31 4</intersection>
<intersection>-22.5 3</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-40.5,62,-40.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-13.5,57.5,-13.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53.5,-22.5,56,-22.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>56,-31,58,-31</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-21.5,65.5,-12.5</points>
<intersection>-21.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-21.5,67.5,-21.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-12.5,65.5,-12.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-32,65.5,-23.5</points>
<intersection>-32 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-32,65.5,-32</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-23.5,67.5,-23.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-41.5,68,-41.5</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>26</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-22.5,73.5,-22.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>N_in0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport>
<gate>
<ID>32</ID>
<type>BE_NOR2</type>
<position>24,-22</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>BE_NOR2</type>
<position>38,-14</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>BE_NOR2</type>
<position>38,-29.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BE_NOR2</type>
<position>48.5,-21.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>BE_NOR2</type>
<position>58.5,-31.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>BE_NOR2</type>
<position>69.5,-40</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>BE_NOR2</type>
<position>80,-31</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>BE_NOR2</type>
<position>69.5,-22.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>BE_NOR2</type>
<position>79.5,-44.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>15.5,-32.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>15.5,-19.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>15.5,-25</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>86,-44.5</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>86,-31</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>24.5,-5.5</position>
<gparam>LABEL_TEXT Full Subtractor Using NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>12,-19</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>12,-24.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>8.5,-32</position>
<gparam>LABEL_TEXT Borrow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>95,-30.5</position>
<gparam>LABEL_TEXT Difference</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>93,-44</position>
<gparam>LABEL_TEXT Borrow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-32.5,55.5,-32.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>55.5 7</intersection>
<intersection>55.5 9</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>55.5,-41,55.5,-32.5</points>
<intersection>-41 8</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>55.5,-41,66.5,-41</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>55.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>55.5,-32.5,55.5,-32.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-21,21,-13</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-19.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-19.5,21,-19.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-13,35,-13</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,-30.5,21,-23</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>-30.5 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-25,21,-25</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>21 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-30.5,35,-30.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>21 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-28.5,31,-15</points>
<intersection>-28.5 3</intersection>
<intersection>-22 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-22,31,-22</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-15,35,-15</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-28.5,35,-28.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-20.5,43,-14</points>
<intersection>-20.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-20.5,45.5,-20.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-14,43,-14</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-45.5,43,-22.5</points>
<intersection>-45.5 3</intersection>
<intersection>-29.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-22.5,45.5,-22.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-29.5,43,-29.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>43,-45.5,76.5,-45.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-30.5,55.5,-21.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-21.5,66.5,-21.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-39,64,-23.5</points>
<intersection>-39 3</intersection>
<intersection>-31.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-23.5,66.5,-23.5</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-31.5,64,-31.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,-39,66.5,-39</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>64 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-43.5,74.5,-32</points>
<intersection>-43.5 3</intersection>
<intersection>-40 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-32,77,-32</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-40,74.5,-40</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>74.5,-43.5,76.5,-43.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-30,74.5,-22.5</points>
<intersection>-30 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-30,77,-30</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-22.5,74.5,-22.5</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-44.5,85,-44.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<connection>
<GID>56</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-31,85,-31</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport>
<gate>
<ID>62</ID>
<type>BA_NAND2</type>
<position>21,-24</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>BA_NAND2</type>
<position>35.5,-15</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>BA_NAND2</type>
<position>35.5,-34</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>BA_NAND2</type>
<position>47.5,-24</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>BA_NAND2</type>
<position>57,-24</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>BA_NAND2</type>
<position>69.5,-15</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_NAND2</type>
<position>68.5,-34.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>BA_NAND2</type>
<position>81.5,-23.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>BA_NAND2</type>
<position>82,-43</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>11,-20.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>11,-28</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>11,-42</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>87.5,-23.5</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>87.5,-43</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>33.5,-4.5</position>
<gparam>LABEL_TEXT Full Subtractor Using NAND gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>7.5,-20</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>7.5,-27.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>10.5,-44</position>
<gparam>LABEL_TEXT Borrow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>97,-23</position>
<gparam>LABEL_TEXT Difference</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>95,-42.5</position>
<gparam>LABEL_TEXT borrow</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-23,18,-14</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-20.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-20.5,18,-20.5</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-14,32.5,-14</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-35,18,-25</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-35 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-28,18,-28</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-35,32.5,-35</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-42,53,-25</points>
<intersection>-42 1</intersection>
<intersection>-35.5 3</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-42,53,-42</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-25,54,-25</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>53,-35.5,65.5,-35.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-44,42.5,-25</points>
<intersection>-44 2</intersection>
<intersection>-34 3</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-25,44.5,-25</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-44,79,-44</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38.5,-34,42.5,-34</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-33,28,-16</points>
<intersection>-33 3</intersection>
<intersection>-24 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-16,32.5,-16</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-24,28,-24</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-33,32.5,-33</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-23,42.5,-15</points>
<intersection>-23 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-23,44.5,-23</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-15,42.5,-15</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-24,52,-23</points>
<intersection>-24 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-23,54,-23</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection>
<intersection>53 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50.5,-24,52,-24</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53,-23,53,-14</points>
<intersection>-23 1</intersection>
<intersection>-14 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>53,-14,66.5,-14</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>53 3</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-33.5,63,-16</points>
<intersection>-33.5 3</intersection>
<intersection>-24 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-16,66.5,-16</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-24,63,-24</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>63,-33.5,65.5,-33.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-22.5,75.5,-15</points>
<intersection>-22.5 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-22.5,78.5,-22.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-15,75.5,-15</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-42,75,-24.5</points>
<intersection>-42 2</intersection>
<intersection>-34.5 1</intersection>
<intersection>-24.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-34.5,75,-34.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-42,79,-42</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>75,-24.5,78.5,-24.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-23.5,86.5,-23.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-43,86.5,-43</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<connection>
<GID>88</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>23,-3.5</position>
<gparam>LABEL_TEXT Full adder using Half adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AI_XOR2</type>
<position>22.5,-16</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AI_XOR2</type>
<position>53.5,-15</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND2</type>
<position>21.5,-30.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND2</type>
<position>52.5,-30.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_OR2</type>
<position>69,-30.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>13,-13.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>13,-19</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>36,-30</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>112</ID>
<type>GA_LED</type>
<position>75,-30.5</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>59.5,-15</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>9.5,-13</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>9.5,-18.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>31.5,-29.5</position>
<gparam>LABEL_TEXT Cin</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>64,-14.5</position>
<gparam>LABEL_TEXT Sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>80,-30</position>
<gparam>LABEL_TEXT Cout</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-35,66,-35</points>
<intersection>24.5 3</intersection>
<intersection>66 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-35,24.5,-30.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>66,-35,66,-31.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-30.5,60.5,-29.5</points>
<intersection>-30.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-29.5,66,-29.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-30.5,60.5,-30.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-29.5,17.5,-13.5</points>
<intersection>-29.5 3</intersection>
<intersection>-15 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-13.5,17.5,-13.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-15,19.5,-15</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>17.5,-29.5,18.5,-29.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-19,19,-17</points>
<intersection>-19 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-19,19,-19</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>16 3</intersection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-17,19.5,-17</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-31.5,16,-19</points>
<intersection>-31.5 4</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,-31.5,18.5,-31.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-16,37.5,-14</points>
<intersection>-16 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-14,50.5,-14</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection>
<intersection>47.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-16,37.5,-16</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,-29.5,47.5,-14</points>
<intersection>-29.5 4</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-29.5,49.5,-29.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>47.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-31.5,43.5,-16</points>
<intersection>-31.5 1</intersection>
<intersection>-30 2</intersection>
<intersection>-16 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-31.5,49.5,-31.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-30,43.5,-30</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-16,50.5,-16</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>72,-30.5,74,-30.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>112</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-15,58.5,-15</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<connection>
<GID>114</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>15.3,-6.425,107.1,-51.8</PageViewport>
<gate>
<ID>194</ID>
<type>AA_TOGGLE</type>
<position>64.5,-14.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>198</ID>
<type>FF_GND</type>
<position>63,-34</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>FF_GND</type>
<position>66,-34</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>GA_LED</type>
<position>54,-40</position>
<input>
<ID>N_in1</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>GA_LED</type>
<position>49.5,-46</position>
<input>
<ID>N_in3</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_TOGGLE</type>
<position>78,-40</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_TOGGLE</type>
<position>70.5,-14.5</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_TOGGLE</type>
<position>72.5,-14.5</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>74.5,-14.5</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_TOGGLE</type>
<position>76.5,-14.5</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>40,-11.5</position>
<gparam>LABEL_TEXT BCD Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_TOGGLE</type>
<position>62.5,-14.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_LABEL</type>
<position>67,-48.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>64.5,-12.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>62.5,-12.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>66.5,-12.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>68.5,-12.5</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>52,-40</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>80.5,-39.5</position>
<gparam>LABEL_TEXT Cin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>65,-48.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>69,-48.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>71,-48.5</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 0.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>158</ID>
<type>AE_FULLADDER_4BIT</type>
<position>68,-41</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>73 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>85 </input>
<input>
<ID>IN_B_0</ID>90 </input>
<input>
<ID>IN_B_1</ID>89 </input>
<input>
<ID>IN_B_2</ID>88 </input>
<input>
<ID>IN_B_3</ID>87 </input>
<output>
<ID>OUT_0</ID>77 </output>
<output>
<ID>OUT_1</ID>76 </output>
<output>
<ID>OUT_2</ID>75 </output>
<output>
<ID>OUT_3</ID>74 </output>
<input>
<ID>carry_in</ID>95 </input>
<output>
<ID>carry_out</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>160</ID>
<type>AE_OR3</type>
<position>41.5,-28.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>56 </input>
<input>
<ID>IN_2</ID>93 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_AND2</type>
<position>55.5,-28.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_AND2</type>
<position>55.5,-33</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_TOGGLE</type>
<position>66.5,-14.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_TOGGLE</type>
<position>68.5,-14.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>65,-46.5</position>
<input>
<ID>N_in3</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>GA_LED</type>
<position>67,-46.5</position>
<input>
<ID>N_in3</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>GA_LED</type>
<position>69,-46.5</position>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>71,-46.5</position>
<input>
<ID>N_in3</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AE_FULLADDER_4BIT</type>
<position>69.5,-23</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>100 </input>
<input>
<ID>IN_B_0</ID>99 </input>
<input>
<ID>IN_B_1</ID>98 </input>
<input>
<ID>IN_B_2</ID>97 </input>
<input>
<ID>IN_B_3</ID>96 </input>
<output>
<ID>OUT_0</ID>90 </output>
<output>
<ID>OUT_1</ID>89 </output>
<output>
<ID>OUT_2</ID>88 </output>
<output>
<ID>OUT_3</ID>87 </output>
<output>
<ID>carry_out</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44.5,-28.5,52.5,-28.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<connection>
<GID>162</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-33,49.5,-30.5</points>
<intersection>-33 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-30.5,49.5,-30.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-33,52.5,-33</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-36,64.5,-36</points>
<intersection>38.5 2</intersection>
<intersection>49.5 6</intersection>
<intersection>64.5 3</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>38.5,-36,38.5,-28.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>64.5,-37,64.5,-36</points>
<intersection>-37 5</intersection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>64,-37,65,-37</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<connection>
<GID>158</GID>
<name>IN_2</name></connection>
<intersection>64.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>49.5,-45,49.5,-36</points>
<connection>
<GID>206</GID>
<name>N_in3</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-45.5,65,-45</points>
<connection>
<GID>178</GID>
<name>N_in3</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-45,66.5,-45</points>
<connection>
<GID>158</GID>
<name>OUT_3</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-45.5,67,-45</points>
<connection>
<GID>180</GID>
<name>N_in3</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-45,67.5,-45</points>
<connection>
<GID>158</GID>
<name>OUT_2</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-45.5,69,-45</points>
<connection>
<GID>182</GID>
<name>N_in3</name></connection>
<intersection>-45 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>68.5,-45,69,-45</points>
<connection>
<GID>158</GID>
<name>OUT_1</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-45.5,71,-45</points>
<connection>
<GID>184</GID>
<name>N_in3</name></connection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-45,71,-45</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-19,66.5,-16.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>-16.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>66.5,-16.5,66.5,-16.5</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-19,68.5,-16.5</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-19 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>67.5,-19,68.5,-19</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-19,65,-16.5</points>
<intersection>-19 3</intersection>
<intersection>-16.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>65,-19,65.5,-19</points>
<intersection>65 0</intersection>
<intersection>65.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>64.5,-16.5,65,-16.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>65.5,-19,65.5,-19</points>
<connection>
<GID>188</GID>
<name>IN_2</name></connection>
<intersection>-19 3</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-37,63,-35</points>
<connection>
<GID>158</GID>
<name>IN_3</name></connection>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-37,66,-35</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-37,70,-32</points>
<connection>
<GID>158</GID>
<name>IN_B_3</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>68,-32,68,-27</points>
<connection>
<GID>188</GID>
<name>OUT_3</name></connection>
<intersection>-32 2</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>68,-32,70,-32</points>
<intersection>68 1</intersection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-27.5,68,-27.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>59 4</intersection>
<intersection>68 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59,-32,59,-27.5</points>
<intersection>-32 6</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>58.5,-32,59,-32</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>59 4</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-37,71,-32</points>
<connection>
<GID>158</GID>
<name>IN_B_2</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>69,-32,69,-27</points>
<connection>
<GID>188</GID>
<name>OUT_2</name></connection>
<intersection>-32 2</intersection>
<intersection>-29.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-32,71,-32</points>
<intersection>69 1</intersection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,-29.5,69,-29.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>69 1</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-37,72,-32</points>
<connection>
<GID>158</GID>
<name>IN_B_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-32,70,-27</points>
<connection>
<GID>188</GID>
<name>OUT_1</name></connection>
<intersection>-32 2</intersection>
<intersection>-31 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70,-32,72,-32</points>
<intersection>70 1</intersection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>59.5,-31,70,-31</points>
<intersection>59.5 4</intersection>
<intersection>70 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59.5,-34,59.5,-31</points>
<intersection>-34 5</intersection>
<intersection>-31 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>58.5,-34,59.5,-34</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>59.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-37,73,-32</points>
<connection>
<GID>158</GID>
<name>IN_B_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>71,-32,71,-27</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>71,-32,73,-32</points>
<intersection>71 1</intersection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-40,60,-40</points>
<connection>
<GID>158</GID>
<name>carry_out</name></connection>
<connection>
<GID>204</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-26.5,49.5,-22</points>
<intersection>-26.5 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-26.5,49.5,-26.5</points>
<connection>
<GID>160</GID>
<name>IN_2</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-22,61.5,-22</points>
<connection>
<GID>188</GID>
<name>carry_out</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-40,76,-40</points>
<connection>
<GID>158</GID>
<name>carry_in</name></connection>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-19,70.5,-16.5</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>-19 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>70.5,-19,71.5,-19</points>
<intersection>70.5 0</intersection>
<intersection>71.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71.5,-19,71.5,-19</points>
<connection>
<GID>188</GID>
<name>IN_B_3</name></connection>
<intersection>-19 4</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>72.5,-19,72.5,-16.5</points>
<connection>
<GID>188</GID>
<name>IN_B_2</name></connection>
<intersection>-16.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>72.5,-16.5,72.5,-16.5</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>72.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>74,-19,74,-16.5</points>
<intersection>-19 3</intersection>
<intersection>-16.5 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>73.5,-19,74,-19</points>
<connection>
<GID>188</GID>
<name>IN_B_1</name></connection>
<intersection>74 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>74,-16.5,74.5,-16.5</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>74 2</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-19,76.5,-16.5</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-19,76.5,-19</points>
<intersection>74.5 2</intersection>
<intersection>76.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>74.5,-19,74.5,-19</points>
<connection>
<GID>188</GID>
<name>IN_B_0</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-19,62.5,-16.5</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-19,64.5,-19</points>
<intersection>62.5 0</intersection>
<intersection>64.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>64.5,-19,64.5,-19</points>
<connection>
<GID>188</GID>
<name>IN_3</name></connection>
<intersection>-19 1</intersection></vsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>